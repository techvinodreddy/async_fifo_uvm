package test_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  
  `include "write_packet.sv"
  `include "write_agent_config.sv"

  `include "read_packet.sv"
  `include "read_agent_config.sv"
  
  `include "environment_config.sv"

  `include "write_sequences.sv"
  `include "write_sequencer.sv"
  `include "write_driver.sv"
  `include "write_monitor.sv"
  `include "write_agent.sv"

  `include "read_sequences.sv"
  `include "read_sequencer.sv"
  `include "read_driver.sv"
  `include "read_monitor.sv"
  `include "read_agent.sv"

  `include "agent_top.sv"

  `include "virtual_sequencer.sv"
  `include "virtual_sequences.sv"
  `include "scoreboard.sv"

  `include "environment.sv"
  `include "test_cases.sv"
endpackage
